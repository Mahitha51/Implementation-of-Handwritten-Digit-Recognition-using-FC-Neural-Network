module fnn_imgclsfctn(input clk,reset,input [27:0] input_image, output nxt_inp,output [3:0] outp)
 

